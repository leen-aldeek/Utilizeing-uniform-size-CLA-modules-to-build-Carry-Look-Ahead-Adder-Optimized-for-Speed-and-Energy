*** SPICE deck for cell 2input_OR{sch} from library IC_Project
*** Created on Fri Jan 10, 2025 16:09:40
*** Last revised on Sat Jan 11, 2025 16:50:20
*** Written on Sat Jan 11, 2025 16:52:43 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: 2input_OR{sch}
Mnmos@0 net@4 A gnd gnd myNMOS L=0.6U W=1.5U
Mnmos@1 net@4 B gnd gnd myNMOS L=0.6U W=1.5U
Mnmos@2 out net@4 gnd gnd myNMOS L=0.6U W=1.5U
Mpmos@0 vdd A net@2 vdd myPMOS L=0.6U W=3U
Mpmos@1 net@2 B net@4 vdd myPMOS L=0.6U W=3U
Mpmos@2 vdd net@4 out vdd myPMOS L=0.6U W=3U

* Spice Code nodes in cell cell '2input_OR{sch}'
* 2-Input OR Gate Implementation
VDD VDD 0 DC 5
VA A 0 PWL 10n 0 20n 5 50n 5 60n 0 70n 0 80n 5 100n 5 110n 0 130n 0 140n 5 170n 5 180n 0 190n 0 200n 5 240n 5 250n 0
VB B 0 PWL 10n 0 20n 5 30n 5 40n 0 50n 0 60n 5 70n 5 80n 0 90n 0 100n 5 110n 5 120n 0 130n 0 140n 5 170n 5 180n 0
* CMOS 2-Input OR Gate
M1 out A 0 0 myNMOS L=0.18u W=1u
M2 out B 0 0 myNMOS L=0.18u W=1u
M3 out A VDD VDD myPMOS L=0.18u W=1u
M4 out B VDD VDD myPMOS L=0.18u W=1u
* Load Capacitance
CLOAD OUT 0 250fF
* Measurement Statements
.measure tran tf TRIG V(out) VAL=4.5 FALL=1 TD=4ns TARG V(OUT) VAL=0.5 FALL=1
.measure tran tr TRIG V(out) VAL=0.5 RISE=1 TD=4ns TARG V(OUT) VAL=4.5 RISE=1
* Transient Analysis
.tran 0 0.5us
* Include Model File
.include "C:\Users\HP\Desktop\electric vlsi\C5_models.txt"
.END
.END
